library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Lab5_Simen_Fuglestad is
	port (
				clk : in std_logic
	);
end entity;

architecture RTL of Lab5_Simen_Fuglestad is
begin
end architecture;